module Not_1 (
input c,
output s);
assign s=!c;
endmodule 