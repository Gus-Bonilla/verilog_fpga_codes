module And_2 (
input a,
input b,
output s);
assign s=a&b;
endmodule 