module Or_2 (
input a,
input b,
output s);
assign s=a|b;
endmodule 