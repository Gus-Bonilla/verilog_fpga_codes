module Mux_2_1 (

input A,
input B,
input C,

output F) ;

//assign F=(~A&C)|(A&B);

//wire W1,W2,W3;		
//
//not (W3,C);
//and (W1,A,W3);
//and (W2,B,C);
//or (F,W1,W2);



endmodule
